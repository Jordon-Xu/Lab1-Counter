module counter #(
    parameter WIDTH = 8
)(
    // interface signals
    input logic              clk,    // clock
    input logic              rst,   // reset
    input logic              en,    // counter enable
    output logic [WIDTH-1:0] count    // clock
);

always_ff @ (posedge clk)
    if (rst) count <= {WIDTH{1'b0}};
    else count <= count + {{WIDTH-1{1'b0}}, en};
        
endmodule

// module counter #(
//     parameter WIDTH = 8
// )(
//     // interface signals
//     input logic clk,       // clock
//     input logic rst,       // reset
//     input logic vbuddy_flag,
//     output logic [WIDTH-1:0] count  // count output
// );

// always_ff @(posedge clk) begin
//     if (rst) begin
//         count <= {WIDTH{1'b0}};
//     end else if (vbuddy_flag) begin 
//         count <= count + {{WIDTH-1{1'b0}},1'b1};
//     end
// end


// endmodule
